module ast

import lexer.token

pub type Statement = LetStatement | ReturnStatement | ExpresionStatement

pub fn (st Statement) token_literal() string {
	return st.token_literal()
}

pub fn (st Statement) str() string {
	return st.str()
}

pub fn (ls LetStatement) token_literal() string {
	return ls.token.value
}

pub fn (ls LetStatement) str() string {
	mut output := ''
	output += '${ls.token_literal()} ${ls.name} = '
	if ls.value != none {
		output += '${ls.value}'
	}
	output += ';'
	return output
}

pub fn (rs ReturnStatement) token_literal() string {
	return rs.token.value
}

pub fn (rs ReturnStatement) str() string {
	mut output := ''
	output += '${rs.token_literal()} '
	if rs.return_value != none {
		output += '${rs.return_value}'
	}
	output += ';'
	return output
}

pub fn (es ExpresionStatement) token_literal() string {
	return es.token.value
}

pub fn (es ExpresionStatement) str() string {
	if es.expression != none {
		return '${es.expression}'
	}
	return ''
}

pub struct ReturnStatement {
pub:
	token        token.TokenType
	return_value ?Expression
}

type Expression = Identifier

pub struct ExpresionStatement {
pub:
	token      token.TokenType
	expression ?Expression
}

pub struct LetStatement {
pub:
	token token.TokenType
	value ?Expression
pub mut:
	name Identifier
}

pub fn (id Identifier) token_literal() string {
	return id.token.value
}

pub fn (id Identifier) str() string {
	return '${id.value}'
}

pub struct Identifier {
pub mut:
	token token.TokenType
	value string
}

pub struct Program {
pub mut:
	statements []Statement
mut:
	idx int
}

fn (mut prog Program) next() ?Statement {
	if prog.idx >= prog.statements.len {
		return none
	}
	defer {
		prog.idx++
	}
	return prog.statements[prog.idx]
}

fn (pro Program) token_literal() string {
	if pro.statements.len > 0 {
		return pro.statements[0].token_literal()
	}
	return ''
}

fn (pro Program) str() string {
	mut output := ''
	return output
}
