module token

pub enum Token {
	assign
	plus
	lparen
	rparen
	lbrace
	rbrace
	comma
	semicolon
	eof
    illegal
}
