module main

struct Items {
	base i32
}

fn main() {
	// data := 'let x = 5 + 5;'
}
