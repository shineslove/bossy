module main

fn main () {

}